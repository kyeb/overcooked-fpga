`timescale 1ns / 1ps

module graphics(
    input reset,
    input clock,
    input [1:0] local_player_ID,
    input [1:0] num_players,
    input logic [2:0] game_state, // welcome screen or 
                  
endmodule
