module action();
endmodule